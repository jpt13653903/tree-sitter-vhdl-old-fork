hello
Hello
HELLO
HeLlO
func
Func
FUNC
FuNc

