func
Func
FUNC
-- A line comment
FuNc
hello
/*
  A multi-line
  block comment
*/
Hello
HELLO
HeLlO
